
package declarations1;

bit [5:0] MAX_QUEUE_SIZE = 'd16;

parameter [7:0] tRC=228;
parameter [7:0] tRAS=152;
parameter [4:0] tRRD_L=22;
parameter [4:0] tRRD_S=14;
parameter [6:0] tRP=76;
parameter [7:0] tRFC=710;
parameter [6:0] tCWD=76;
parameter [6:0] tCL=80;
parameter [6:0] tRCD=76;
parameter [5:0] tWR=60;
parameter [5:0] tRTP=36;
parameter [4:0] tCCD_L=22;
parameter [4:0] tCCD_S=14;
parameter [6:0] tCCD_L_WR=94;
parameter [4:0] tCCD_S_WR=14;
parameter [4:0] tBURST=16;
parameter [5:0] tCCD_L_RTW=30;
parameter [5:0] tCCD_S_RTW=30;
parameter [7:0] tCCD_L_WTR=138;
parameter [6:0] tCCD_S_WTR=102;

endpackage