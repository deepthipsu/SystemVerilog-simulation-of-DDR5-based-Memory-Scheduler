
module test;



endmodule