
package declarations1;

bit[5:0] MAX_QUEUE_SIZE = 'd16;

endpackage